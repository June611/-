module aenum();
enum {s[5]} state;

initial begin
state =s4;
state =s5;
end
endmodule
