module FSM();
	enum{GO, STOP} fsm1_state;
	enum{GO, WAIT,DONE} fsm2_state;	//GO already have a value

endmodule