package chip_types;
    typedef enum {FETCH, WRITE, ADD, SUB, MULT, DIV, SHIFT, NOP} instr_t;
endpackage

import chip_types::*;

module controller(output logic read, write,
                    input instr_t instruction,
                    input wire clk, resetN );
    enum {WAIT, LOAD, STORE} state, nextState;

   always @(posedge clk, negedge resetN)
        if(!resetN) state = WAIT;
        else state = nextState;

    always @(state) begin
        case(state)
            WAIT:nextState = LOAD;
            LOAD:nextState = STORE;
            STORE: nextState = WAIT;
        endcase
    end

    always@(state, instruction)begin
        read = 0; write=0;
        if(state == LOAD && instruction ==FETCH)    read = 1;
        else if(state == STORE && instruction == WRITE) write=1;
    end

	initial begin
		#5 state = WAIT;
		#5 instruction = FETCH;
		//#10 state = LOAD;
	end
endmodule
