module aenum();
enum {s[5]} state;

initial
state =s5;

endmodule
