module compressed_array();

	bit [31:0] a;
	logic [4:0]b;
	byte [7:0] c;
endmodule