module test();
	enum logic {ON = 1'b0, OFF = 1'b1, HI = 1'bz, UN = 1'bx} four_st;

endmodule